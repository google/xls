// Copyright 2021 The XLS Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module isqrt(num, out);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  (* src = "/tmp/sqrt.cc.v:2.21-2.24" *)
  input [15:0] num;
  (* src = "/tmp/sqrt.cc.v:3.21-3.24" *)
  output [7:0] out;
  inv _197_ (
    .A(num[15]),
    .Y(_126_)
  );
  inv _198_ (
    .A(num[12]),
    .Y(_127_)
  );
  inv _199_ (
    .A(num[8]),
    .Y(_128_)
  );
  inv _200_ (
    .A(num[9]),
    .Y(_129_)
  );
  inv _201_ (
    .A(num[10]),
    .Y(_130_)
  );
  inv _202_ (
    .A(num[4]),
    .Y(_131_)
  );
  inv _203_ (
    .A(num[5]),
    .Y(_132_)
  );
  inv _204_ (
    .A(num[6]),
    .Y(_133_)
  );
  inv _205_ (
    .A(num[7]),
    .Y(_134_)
  );
  inv _206_ (
    .A(num[3]),
    .Y(_135_)
  );
  inv _207_ (
    .A(num[2]),
    .Y(_136_)
  );
  orny2 _208_ (
    .A(num[14]),
    .B(num[15]),
    .Y(_137_)
  );
  inv _209_ (
    .A(_137_),
    .Y(out[7])
  );
  nor2 _210_ (
    .A(num[15]),
    .B(num[14]),
    .Y(_138_)
  );
  or2 _211_ (
    .A(num[12]),
    .B(num[13]),
    .Y(_139_)
  );
  nand2 _212_ (
    .A(_138_),
    .B(_139_),
    .Y(_140_)
  );
  inv _213_ (
    .A(_140_),
    .Y(out[6])
  );
  nand2 _214_ (
    .A(_127_),
    .B(_138_),
    .Y(_141_)
  );
  and2 _215_ (
    .A(num[13]),
    .B(_141_),
    .Y(_142_)
  );
  nand2 _216_ (
    .A(_137_),
    .B(_142_),
    .Y(_143_)
  );
  or2 _217_ (
    .A(num[10]),
    .B(num[11]),
    .Y(_144_)
  );
  or2 _218_ (
    .A(num[13]),
    .B(_137_),
    .Y(_145_)
  );
  and2 _219_ (
    .A(_144_),
    .B(_145_),
    .Y(_146_)
  );
  nand2 _220_ (
    .A(_143_),
    .B(_146_),
    .Y(_147_)
  );
  nand2 _221_ (
    .A(_127_),
    .B(_147_),
    .Y(_148_)
  );
  and2 _222_ (
    .A(_126_),
    .B(_148_),
    .Y(_149_)
  );
  orny2 _223_ (
    .A(num[12]),
    .B(num[13]),
    .Y(_150_)
  );
  nand2 _224_ (
    .A(_149_),
    .B(_150_),
    .Y(_151_)
  );
  inv _225_ (
    .A(_151_),
    .Y(out[5])
  );
  andny2 _226_ (
    .A(_151_),
    .B(_130_),
    .Y(_152_)
  );
  imux2 _227_ (
    .A(_140_),
    .B(_144_),
    .S(_151_),
    .Y(_153_)
  );
  xnor2 _228_ (
    .A(num[12]),
    .B(_153_),
    .Y(_154_)
  );
  nand2 _229_ (
    .A(_137_),
    .B(_154_),
    .Y(_155_)
  );
  xnor2 _230_ (
    .A(out[7]),
    .B(_154_),
    .Y(_156_)
  );
  xnor2 _231_ (
    .A(num[11]),
    .B(_152_),
    .Y(_157_)
  );
  inv _232_ (
    .A(_157_),
    .Y(_158_)
  );
  or2 _233_ (
    .A(out[6]),
    .B(_157_),
    .Y(_159_)
  );
  xnor2 _234_ (
    .A(_140_),
    .B(_157_),
    .Y(_160_)
  );
  nor2 _235_ (
    .A(num[8]),
    .B(num[9]),
    .Y(_161_)
  );
  imux2 _236_ (
    .A(out[5]),
    .B(_161_),
    .S(num[10]),
    .Y(_162_)
  );
  inv _237_ (
    .A(_162_),
    .Y(_163_)
  );
  nand2 _238_ (
    .A(_160_),
    .B(_163_),
    .Y(_164_)
  );
  nand2 _239_ (
    .A(_159_),
    .B(_164_),
    .Y(_165_)
  );
  nand2 _240_ (
    .A(_156_),
    .B(_165_),
    .Y(_166_)
  );
  orny2 _241_ (
    .A(_142_),
    .B(_149_),
    .Y(_167_)
  );
  and2 _242_ (
    .A(_155_),
    .B(_167_),
    .Y(_168_)
  );
  nand2 _243_ (
    .A(_166_),
    .B(_168_),
    .Y(_169_)
  );
  nand2 _244_ (
    .A(_126_),
    .B(_169_),
    .Y(_170_)
  );
  inv _245_ (
    .A(_170_),
    .Y(out[4])
  );
  xnor2 _246_ (
    .A(_160_),
    .B(_162_),
    .Y(_171_)
  );
  imux2 _247_ (
    .A(_158_),
    .B(_171_),
    .S(_170_),
    .Y(_172_)
  );
  nand2 _248_ (
    .A(_137_),
    .B(_172_),
    .Y(_173_)
  );
  xnor2 _249_ (
    .A(out[7]),
    .B(_172_),
    .Y(_174_)
  );
  xnor2 _250_ (
    .A(_130_),
    .B(_151_),
    .Y(_175_)
  );
  xnor2 _251_ (
    .A(num[10]),
    .B(_161_),
    .Y(_176_)
  );
  imux2 _252_ (
    .A(_175_),
    .B(_176_),
    .S(_170_),
    .Y(_177_)
  );
  or2 _253_ (
    .A(out[6]),
    .B(_177_),
    .Y(_178_)
  );
  xnor2 _254_ (
    .A(out[6]),
    .B(_177_),
    .Y(_179_)
  );
  andny2 _255_ (
    .A(_170_),
    .B(_128_),
    .Y(_180_)
  );
  xnor2 _256_ (
    .A(_129_),
    .B(_180_),
    .Y(_181_)
  );
  nand2 _257_ (
    .A(_151_),
    .B(_181_),
    .Y(_182_)
  );
  xnor2 _258_ (
    .A(out[5]),
    .B(_181_),
    .Y(_183_)
  );
  nor2 _259_ (
    .A(num[6]),
    .B(num[7]),
    .Y(_184_)
  );
  imux2 _260_ (
    .A(out[4]),
    .B(_184_),
    .S(num[8]),
    .Y(_185_)
  );
  inv _261_ (
    .A(_185_),
    .Y(_186_)
  );
  nand2 _262_ (
    .A(_183_),
    .B(_186_),
    .Y(_187_)
  );
  and2 _263_ (
    .A(_182_),
    .B(_187_),
    .Y(_188_)
  );
  or2 _264_ (
    .A(_179_),
    .B(_188_),
    .Y(_189_)
  );
  nand2 _265_ (
    .A(_178_),
    .B(_189_),
    .Y(_190_)
  );
  nand2 _266_ (
    .A(_174_),
    .B(_190_),
    .Y(_191_)
  );
  xor2 _267_ (
    .A(_156_),
    .B(_165_),
    .Y(_192_)
  );
  andny2 _268_ (
    .A(_170_),
    .B(_192_),
    .Y(_193_)
  );
  orny2 _269_ (
    .A(_154_),
    .B(_169_),
    .Y(_194_)
  );
  andny2 _270_ (
    .A(_193_),
    .B(_194_),
    .Y(_195_)
  );
  and2 _271_ (
    .A(_173_),
    .B(_195_),
    .Y(_196_)
  );
  nand2 _272_ (
    .A(_191_),
    .B(_196_),
    .Y(_000_)
  );
  nand2 _273_ (
    .A(_126_),
    .B(_000_),
    .Y(_001_)
  );
  inv _274_ (
    .A(_001_),
    .Y(out[3])
  );
  xnor2 _275_ (
    .A(_179_),
    .B(_188_),
    .Y(_002_)
  );
  imux2 _276_ (
    .A(_177_),
    .B(_002_),
    .S(_001_),
    .Y(_003_)
  );
  or2 _277_ (
    .A(out[7]),
    .B(_003_),
    .Y(_004_)
  );
  xnor2 _278_ (
    .A(_137_),
    .B(_003_),
    .Y(_005_)
  );
  xnor2 _279_ (
    .A(_183_),
    .B(_185_),
    .Y(_006_)
  );
  imux2 _280_ (
    .A(_181_),
    .B(_006_),
    .S(_001_),
    .Y(_007_)
  );
  inv _281_ (
    .A(_007_),
    .Y(_008_)
  );
  nand2 _282_ (
    .A(_140_),
    .B(_007_),
    .Y(_009_)
  );
  xnor2 _283_ (
    .A(_140_),
    .B(_007_),
    .Y(_010_)
  );
  xnor2 _284_ (
    .A(_128_),
    .B(_170_),
    .Y(_011_)
  );
  xnor2 _285_ (
    .A(num[8]),
    .B(_184_),
    .Y(_012_)
  );
  imux2 _286_ (
    .A(_011_),
    .B(_012_),
    .S(_001_),
    .Y(_013_)
  );
  or2 _287_ (
    .A(out[5]),
    .B(_013_),
    .Y(_014_)
  );
  andny2 _288_ (
    .A(_001_),
    .B(_133_),
    .Y(_015_)
  );
  xnor2 _289_ (
    .A(_134_),
    .B(_015_),
    .Y(_016_)
  );
  inv _290_ (
    .A(_016_),
    .Y(_017_)
  );
  nand2 _291_ (
    .A(_170_),
    .B(_016_),
    .Y(_018_)
  );
  xnor2 _292_ (
    .A(out[4]),
    .B(_016_),
    .Y(_019_)
  );
  nor2 _293_ (
    .A(num[4]),
    .B(num[5]),
    .Y(_020_)
  );
  imux2 _294_ (
    .A(out[3]),
    .B(_020_),
    .S(num[6]),
    .Y(_021_)
  );
  inv _295_ (
    .A(_021_),
    .Y(_022_)
  );
  nand2 _296_ (
    .A(_019_),
    .B(_022_),
    .Y(_023_)
  );
  nand2 _297_ (
    .A(_018_),
    .B(_023_),
    .Y(_024_)
  );
  xnor2 _298_ (
    .A(_151_),
    .B(_013_),
    .Y(_025_)
  );
  nand2 _299_ (
    .A(_024_),
    .B(_025_),
    .Y(_026_)
  );
  and2 _300_ (
    .A(_014_),
    .B(_026_),
    .Y(_027_)
  );
  or2 _301_ (
    .A(_010_),
    .B(_027_),
    .Y(_028_)
  );
  nand2 _302_ (
    .A(_009_),
    .B(_028_),
    .Y(_029_)
  );
  nand2 _303_ (
    .A(_005_),
    .B(_029_),
    .Y(_030_)
  );
  xor2 _304_ (
    .A(_174_),
    .B(_190_),
    .Y(_031_)
  );
  imux2 _305_ (
    .A(_172_),
    .B(_031_),
    .S(_001_),
    .Y(_032_)
  );
  andyn2 _306_ (
    .A(_004_),
    .B(_032_),
    .Y(_033_)
  );
  nand2 _307_ (
    .A(_030_),
    .B(_033_),
    .Y(_034_)
  );
  nand2 _308_ (
    .A(_126_),
    .B(_034_),
    .Y(_035_)
  );
  inv _309_ (
    .A(_035_),
    .Y(out[2])
  );
  xnor2 _310_ (
    .A(_024_),
    .B(_025_),
    .Y(_036_)
  );
  imux2 _311_ (
    .A(_013_),
    .B(_036_),
    .S(_035_),
    .Y(_037_)
  );
  inv _312_ (
    .A(_037_),
    .Y(_038_)
  );
  or2 _313_ (
    .A(out[6]),
    .B(_037_),
    .Y(_039_)
  );
  xnor2 _314_ (
    .A(_140_),
    .B(_037_),
    .Y(_040_)
  );
  inv _315_ (
    .A(_040_),
    .Y(_041_)
  );
  xnor2 _316_ (
    .A(_019_),
    .B(_022_),
    .Y(_042_)
  );
  imux2 _317_ (
    .A(_017_),
    .B(_042_),
    .S(_035_),
    .Y(_043_)
  );
  inv _318_ (
    .A(_043_),
    .Y(_044_)
  );
  or2 _319_ (
    .A(out[5]),
    .B(_043_),
    .Y(_045_)
  );
  xnor2 _320_ (
    .A(_151_),
    .B(_043_),
    .Y(_046_)
  );
  inv _321_ (
    .A(_046_),
    .Y(_047_)
  );
  xnor2 _322_ (
    .A(_133_),
    .B(_001_),
    .Y(_048_)
  );
  xnor2 _323_ (
    .A(num[6]),
    .B(_020_),
    .Y(_049_)
  );
  imux2 _324_ (
    .A(_048_),
    .B(_049_),
    .S(_035_),
    .Y(_050_)
  );
  inv _325_ (
    .A(_050_),
    .Y(_051_)
  );
  or2 _326_ (
    .A(out[4]),
    .B(_050_),
    .Y(_052_)
  );
  xnor2 _327_ (
    .A(_170_),
    .B(_050_),
    .Y(_053_)
  );
  inv _328_ (
    .A(_053_),
    .Y(_054_)
  );
  andny2 _329_ (
    .A(_035_),
    .B(_131_),
    .Y(_055_)
  );
  xnor2 _330_ (
    .A(_132_),
    .B(_055_),
    .Y(_056_)
  );
  nand2 _331_ (
    .A(_001_),
    .B(_056_),
    .Y(_057_)
  );
  xnor2 _332_ (
    .A(out[3]),
    .B(_056_),
    .Y(_058_)
  );
  nor2 _333_ (
    .A(num[3]),
    .B(num[2]),
    .Y(_059_)
  );
  imux2 _334_ (
    .A(out[2]),
    .B(_059_),
    .S(num[4]),
    .Y(_060_)
  );
  inv _335_ (
    .A(_060_),
    .Y(_061_)
  );
  nand2 _336_ (
    .A(_058_),
    .B(_061_),
    .Y(_062_)
  );
  and2 _337_ (
    .A(_057_),
    .B(_062_),
    .Y(_063_)
  );
  or2 _338_ (
    .A(_054_),
    .B(_063_),
    .Y(_064_)
  );
  and2 _339_ (
    .A(_052_),
    .B(_064_),
    .Y(_065_)
  );
  or2 _340_ (
    .A(_047_),
    .B(_065_),
    .Y(_066_)
  );
  and2 _341_ (
    .A(_045_),
    .B(_066_),
    .Y(_067_)
  );
  or2 _342_ (
    .A(_041_),
    .B(_067_),
    .Y(_068_)
  );
  nand2 _343_ (
    .A(_039_),
    .B(_068_),
    .Y(_069_)
  );
  xnor2 _344_ (
    .A(_010_),
    .B(_027_),
    .Y(_070_)
  );
  imux2 _345_ (
    .A(_008_),
    .B(_070_),
    .S(_035_),
    .Y(_071_)
  );
  or2 _346_ (
    .A(out[7]),
    .B(_071_),
    .Y(_072_)
  );
  xnor2 _347_ (
    .A(_137_),
    .B(_071_),
    .Y(_073_)
  );
  nand2 _348_ (
    .A(_069_),
    .B(_073_),
    .Y(_074_)
  );
  xnor2 _349_ (
    .A(_005_),
    .B(_029_),
    .Y(_075_)
  );
  imux2 _350_ (
    .A(_003_),
    .B(_075_),
    .S(_035_),
    .Y(_076_)
  );
  and2 _351_ (
    .A(_072_),
    .B(_076_),
    .Y(_077_)
  );
  nand2 _352_ (
    .A(_074_),
    .B(_077_),
    .Y(_078_)
  );
  nand2 _353_ (
    .A(_126_),
    .B(_078_),
    .Y(_079_)
  );
  inv _354_ (
    .A(_079_),
    .Y(out[1])
  );
  xnor2 _355_ (
    .A(_040_),
    .B(_067_),
    .Y(_080_)
  );
  imux2 _356_ (
    .A(_038_),
    .B(_080_),
    .S(_079_),
    .Y(_081_)
  );
  or2 _357_ (
    .A(_137_),
    .B(_081_),
    .Y(_082_)
  );
  xnor2 _358_ (
    .A(_046_),
    .B(_065_),
    .Y(_083_)
  );
  imux2 _359_ (
    .A(_044_),
    .B(_083_),
    .S(_079_),
    .Y(_084_)
  );
  nand2 _360_ (
    .A(_140_),
    .B(_084_),
    .Y(_085_)
  );
  xnor2 _361_ (
    .A(num[4]),
    .B(_035_),
    .Y(_086_)
  );
  xnor2 _362_ (
    .A(_131_),
    .B(_059_),
    .Y(_087_)
  );
  imux2 _363_ (
    .A(_086_),
    .B(_087_),
    .S(_079_),
    .Y(_088_)
  );
  nand2 _364_ (
    .A(_001_),
    .B(_088_),
    .Y(_089_)
  );
  nor2 _365_ (
    .A(num[0]),
    .B(num[1]),
    .Y(_090_)
  );
  nand2 _366_ (
    .A(_136_),
    .B(_090_),
    .Y(_091_)
  );
  nand2 _367_ (
    .A(_035_),
    .B(_091_),
    .Y(_092_)
  );
  xnor2 _368_ (
    .A(_135_),
    .B(_079_),
    .Y(_093_)
  );
  nand2 _369_ (
    .A(_092_),
    .B(_093_),
    .Y(_094_)
  );
  or2 _370_ (
    .A(_035_),
    .B(_091_),
    .Y(_095_)
  );
  andny2 _371_ (
    .A(num[3]),
    .B(num[2]),
    .Y(_096_)
  );
  andny2 _372_ (
    .A(_079_),
    .B(_096_),
    .Y(_097_)
  );
  andyn2 _373_ (
    .A(_095_),
    .B(_097_),
    .Y(_098_)
  );
  nand2 _374_ (
    .A(_094_),
    .B(_098_),
    .Y(_099_)
  );
  nand2 _375_ (
    .A(_089_),
    .B(_099_),
    .Y(_100_)
  );
  xnor2 _376_ (
    .A(_058_),
    .B(_060_),
    .Y(_101_)
  );
  imux2 _377_ (
    .A(_056_),
    .B(_101_),
    .S(_079_),
    .Y(_102_)
  );
  or2 _378_ (
    .A(_170_),
    .B(_102_),
    .Y(_103_)
  );
  or2 _379_ (
    .A(_001_),
    .B(_088_),
    .Y(_104_)
  );
  and2 _380_ (
    .A(_103_),
    .B(_104_),
    .Y(_105_)
  );
  nand2 _381_ (
    .A(_100_),
    .B(_105_),
    .Y(_106_)
  );
  xnor2 _382_ (
    .A(_053_),
    .B(_063_),
    .Y(_107_)
  );
  imux2 _383_ (
    .A(_051_),
    .B(_107_),
    .S(_079_),
    .Y(_108_)
  );
  nand2 _384_ (
    .A(_151_),
    .B(_108_),
    .Y(_109_)
  );
  nand2 _385_ (
    .A(_170_),
    .B(_102_),
    .Y(_110_)
  );
  and2 _386_ (
    .A(_109_),
    .B(_110_),
    .Y(_111_)
  );
  nand2 _387_ (
    .A(_106_),
    .B(_111_),
    .Y(_112_)
  );
  or2 _388_ (
    .A(_140_),
    .B(_084_),
    .Y(_113_)
  );
  or2 _389_ (
    .A(_151_),
    .B(_108_),
    .Y(_114_)
  );
  and2 _390_ (
    .A(_113_),
    .B(_114_),
    .Y(_115_)
  );
  nand2 _391_ (
    .A(_112_),
    .B(_115_),
    .Y(_116_)
  );
  nand2 _392_ (
    .A(_085_),
    .B(_116_),
    .Y(_117_)
  );
  nand2 _393_ (
    .A(_082_),
    .B(_117_),
    .Y(_118_)
  );
  nand2 _394_ (
    .A(_137_),
    .B(_081_),
    .Y(_119_)
  );
  xnor2 _395_ (
    .A(_069_),
    .B(_073_),
    .Y(_120_)
  );
  and2 _396_ (
    .A(_071_),
    .B(_076_),
    .Y(_121_)
  );
  and2 _397_ (
    .A(_126_),
    .B(_121_),
    .Y(_122_)
  );
  imux2 _398_ (
    .A(_122_),
    .B(_120_),
    .S(_079_),
    .Y(_123_)
  );
  and2 _399_ (
    .A(_119_),
    .B(_123_),
    .Y(_124_)
  );
  nand2 _400_ (
    .A(_118_),
    .B(_124_),
    .Y(_125_)
  );
  and2 _401_ (
    .A(_126_),
    .B(_125_),
    .Y(out[0])
  );
endmodule
