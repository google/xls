module __axi_reader__AxiReaderInternalRInst__AxiReaderInternalR_0__16_128_16_8_8_5_4_12_next(
  input wire clk,
  input wire rst,
  input wire [139:0] axi_reader__axi_r_r_data,
  input wire axi_reader__axi_r_r_vld,
  input wire axi_reader__axi_st_s_rdy,
  input wire [47:0] axi_reader__conf_r_data,
  input wire axi_reader__conf_r_vld,
  input wire axi_reader__resp_s_rdy,
  output wire axi_reader__axi_r_r_rdy,
  output wire [176:0] axi_reader__axi_st_s_data,
  output wire axi_reader__axi_st_s_vld,
  output wire axi_reader__conf_r_rdy,
  output wire axi_reader__resp_s_data,
  output wire axi_reader__resp_s_vld
);
  wire [47:0] __axi_reader__conf_r_data_reg_init = {16'h0000, 16'h0000, 8'h00, 4'h0, 4'h0};
  wire [47:0] __axi_reader__conf_r_data_skid_reg_init = {16'h0000, 16'h0000, 8'h00, 4'h0, 4'h0};
  wire [139:0] __axi_reader__axi_r_r_data_reg_init = {8'h00, 128'h0000_0000_0000_0000_0000_0000_0000_0000, 3'h0, 1'h0};
  wire [139:0] __axi_reader__axi_r_r_data_skid_reg_init = {8'h00, 128'h0000_0000_0000_0000_0000_0000_0000_0000, 3'h0, 1'h0};
  wire [176:0] __axi_reader__axi_st_s_data_reg_init = {128'h0000_0000_0000_0000_0000_0000_0000_0000, 16'h0000, 16'h0000, 8'h00, 8'h00, 1'h0};
  wire [176:0] __axi_reader__axi_st_s_data_skid_reg_init = {128'h0000_0000_0000_0000_0000_0000_0000_0000, 16'h0000, 16'h0000, 8'h00, 8'h00, 1'h0};
  wire [139:0] literal_2163 = {8'h00, 128'h0000_0000_0000_0000_0000_0000_0000_0000, 3'h0, 1'h0};
  wire [47:0] literal_1942 = {16'h0000, 16'h0000, 8'h00, 4'h0, 4'h0};
  reg [3:0] ____state_4;
  reg [3:0] ____state_5;
  reg [7:0] ____state_3;
  reg ____state_0;
  reg [15:0] ____state_2;
  reg p0_____state_0__1;
  reg [3:0] p0_____state_4__1;
  reg [3:0] p0_____state_5__1;
  reg p0_eq_1885;
  reg [5:0] p0_sel_1917;
  reg p0_ugt_1918;
  reg p0_eq_1928;
  reg p0_not_1927;
  reg p0_and_1940;
  reg p0_and_1929;
  reg p1_____state_0__1;
  reg [10:0] p1_sel_2098;
  reg p1_ugt_2102;
  reg p1_ugt_2110;
  reg p1_ugt_2118;
  reg p1_eq_1928;
  reg [15:0] p1_and_2124;
  reg p1_not_1927;
  reg p1_and_1940;
  reg p1_and_1929;
  reg p0_valid;
  reg p1_valid;
  reg __axi_reader__axi_st_s_data_has_been_sent_reg;
  reg __axi_reader__resp_s_data_has_been_sent_reg;
  reg [47:0] __axi_reader__conf_r_data_reg;
  reg [47:0] __axi_reader__conf_r_data_skid_reg;
  reg __axi_reader__conf_r_data_valid_reg;
  reg __axi_reader__conf_r_data_valid_skid_reg;
  reg [139:0] __axi_reader__axi_r_r_data_reg;
  reg [139:0] __axi_reader__axi_r_r_data_skid_reg;
  reg __axi_reader__axi_r_r_data_valid_reg;
  reg __axi_reader__axi_r_r_data_valid_skid_reg;
  reg [176:0] __axi_reader__axi_st_s_data_reg;
  reg [176:0] __axi_reader__axi_st_s_data_skid_reg;
  reg __axi_reader__axi_st_s_data_valid_reg;
  reg __axi_reader__axi_st_s_data_valid_skid_reg;
  reg __axi_reader__resp_s_data_reg;
  reg __axi_reader__resp_s_data_skid_reg;
  reg __axi_reader__resp_s_data_valid_reg;
  reg __axi_reader__resp_s_data_valid_skid_reg;
  wire [15:0] and_2019;
  wire [15:0] and_2031;
  wire [15:0] and_2047;
  wire [139:0] axi_reader__axi_r_r_data_select;
  wire [139:0] axi_reader__axi_r_r_select;
  wire [2:0] axi_r_resp;
  wire is_err;
  wire [15:0] and_2070;
  wire nor_2181;
  wire axi_reader__axi_st_s_not_pred;
  wire axi_reader__axi_st_s_data_from_skid_rdy;
  wire axi_reader__resp_s_data_from_skid_rdy;
  wire or_2416;
  wire p2_all_active_outputs_ready;
  wire [15:0] and_2094;
  wire p2_stage_done;
  wire p2_not_valid;
  wire is_last_group;
  wire not_1927;
  wire p1_enable;
  wire and_1929;
  wire nor_1930;
  wire [2:0] sel_1900;
  wire p1_data_enable;
  wire p1_not_valid;
  wire [13:0] concat_2156;
  wire [1:0] ____state_2__next_value_predicates;
  wire [2:0] ____state_3__next_value_predicates;
  wire [1:0] ____state_4__next_value_predicates;
  wire [8:0] concat_2068;
  wire [3:0] MAX_LANE__2;
  wire p0_enable;
  wire p0_stage_done;
  wire [2:0] one_hot_1937;
  wire [3:0] one_hot_1938;
  wire [2:0] one_hot_1939;
  wire [15:0] and_2111;
  wire p0_data_enable;
  wire __axi_reader__axi_st_s_vld_buf;
  wire __axi_reader__axi_st_s_data_not_has_been_sent;
  wire __axi_reader__resp_s_vld_buf;
  wire __axi_reader__resp_s_data_not_has_been_sent;
  wire [47:0] axi_reader__conf_r_data_select;
  wire axi_reader__conf_r_data_from_skid_rdy;
  wire and_2270;
  wire axi_reader__axi_r_r_data_from_skid_rdy;
  wire and_2271;
  wire [14:0] high_mask_squeezed;
  wire high_mask_squeezed_const_lsb_bits;
  wire __axi_reader__axi_st_s_data_valid_and_not_has_been_sent;
  wire __axi_reader__resp_s_data_valid_and_not_has_been_sent;
  wire [3:0] MAX_LANE;
  wire and_2242;
  wire [47:0] axi_reader__conf_r_select;
  wire and_2249;
  wire and_2256;
  wire axi_reader__conf_r_data_data_valid_load_en;
  wire axi_reader__conf_r_data_to_is_not_rdy;
  wire axi_reader__axi_r_r_data_data_valid_load_en;
  wire axi_reader__axi_r_r_data_to_is_not_rdy;
  wire [15:0] low_mask;
  wire [15:0] high_mask;
  wire axi_reader__axi_st_s_data_data_valid_load_en;
  wire axi_reader__axi_st_s_data_to_is_not_rdy;
  wire axi_reader__resp_s_data_data_valid_load_en;
  wire axi_reader__resp_s_data_to_is_not_rdy;
  wire ____state_2__at_most_one_next_value;
  wire ____state_3__at_most_one_next_value;
  wire ____state_4__at_most_one_next_value;
  wire [10:0] concat_2092;
  wire [5:0] concat_1914;
  wire [3:0] high_lane;
  wire [3:0] MAX_LANE__1;
  wire is_last_tran;
  wire [1:0] concat_2244;
  wire [2:0] concat_2251;
  wire [7:0] add_1968;
  wire [1:0] concat_2257;
  wire __axi_reader__axi_st_s_data_valid_and_all_active_outputs_ready;
  wire __axi_reader__resp_s_data_valid_and_all_active_outputs_ready;
  wire axi_reader__conf_r_data_data_is_sent_to;
  wire axi_reader__conf_r_data_skid_data_load_en;
  wire axi_reader__conf_r_data_skid_valid_set_zero;
  wire axi_reader__axi_r_r_data_data_is_sent_to;
  wire axi_reader__axi_r_r_data_skid_data_load_en;
  wire axi_reader__axi_r_r_data_skid_valid_set_zero;
  wire [127:0] axi_r_data;
  wire [15:0] mask;
  wire axi_reader__axi_st_s_data_data_is_sent_to;
  wire axi_reader__axi_st_s_data_skid_data_load_en;
  wire axi_reader__axi_st_s_data_skid_valid_set_zero;
  wire axi_reader__resp_s_data_data_is_sent_to;
  wire axi_reader__resp_s_data_skid_data_load_en;
  wire axi_reader__resp_s_data_skid_valid_set_zero;
  wire [176:0] axi_reader__axi_st_s_data_select;
  wire axi_reader__axi_st_s_data_valid_or;
  wire axi_reader__resp_s_data_select;
  wire axi_reader__resp_s_data_valid_or;
  wire or_2408;
  wire [10:0] sel_2098;
  wire ugt_2102;
  wire ugt_2110;
  wire ugt_2118;
  wire [15:0] and_2124;
  wire eq_1885;
  wire [5:0] sel_1917;
  wire ugt_1918;
  wire eq_1928;
  wire and_1940;
  wire nand_1961;
  wire [15:0] one_hot_sel_2245;
  wire or_2246;
  wire [7:0] one_hot_sel_2252;
  wire or_2253;
  wire [3:0] one_hot_sel_2258;
  wire or_2259;
  wire [3:0] one_hot_sel_2265;
  wire __axi_reader__axi_st_s_data_not_stage_load;
  wire __axi_reader__axi_st_s_data_has_been_sent_reg_load_en;
  wire __axi_reader__resp_s_data_not_stage_load;
  wire __axi_reader__resp_s_data_has_been_sent_reg_load_en;
  wire axi_reader__conf_r_data_data_valid_load_en__1;
  wire axi_reader__conf_r_data_skid_valid_load_en;
  wire axi_reader__axi_r_r_data_data_valid_load_en__1;
  wire axi_reader__axi_r_r_data_skid_valid_load_en;
  wire [176:0] __axi_reader__axi_st_s_data_buf;
  wire axi_reader__axi_st_s_data_data_valid_load_en__1;
  wire axi_reader__axi_st_s_data_skid_valid_load_en;
  wire axi_reader__resp_s_data_data_valid_load_en__1;
  wire axi_reader__resp_s_data_skid_valid_load_en;
  assign and_2019 = ({15'h0001, ~p0_____state_4__1[0]} & {16{p0_eq_1885}} | 16'h0004) & {16{~(&p0_____state_4__1[1:0])}};
  assign and_2031 = ((and_2019 | 16'h0008) & {16{~p0_____state_4__1[2]}} | 16'h0010) & {16{p0_____state_4__1 < 4'h5}};
  assign and_2047 = ((and_2031 | 16'h0020) & {16{p0_____state_4__1 < 4'h6}} | 16'h0040) & {16{~(&p0_____state_4__1[2:0])}};
  assign axi_reader__axi_r_r_data_select = __axi_reader__axi_r_r_data_valid_skid_reg ? __axi_reader__axi_r_r_data_skid_reg : __axi_reader__axi_r_r_data_reg;
  assign axi_reader__axi_r_r_select = p1_____state_0__1 ? axi_reader__axi_r_r_data_select : literal_2163;
  assign axi_r_resp = axi_reader__axi_r_r_select[3:1];
  assign is_err = axi_r_resp != 3'h0;
  assign and_2070 = ((and_2047 | 16'h0080) & {16{~p0_____state_4__1[3]}} | 16'h0100) & {16{p0_____state_4__1 < 4'h9}};
  assign nor_2181 = ~(p1_not_1927 | is_err);
  assign axi_reader__axi_st_s_not_pred = ~nor_2181;
  assign axi_reader__axi_st_s_data_from_skid_rdy = ~__axi_reader__axi_st_s_data_valid_skid_reg;
  assign axi_reader__resp_s_data_from_skid_rdy = ~__axi_reader__resp_s_data_valid_skid_reg;
  assign or_2416 = ~p1_____state_0__1 | __axi_reader__axi_r_r_data_valid_reg | __axi_reader__axi_r_r_data_valid_skid_reg;
  assign p2_all_active_outputs_ready = (axi_reader__axi_st_s_not_pred | axi_reader__axi_st_s_data_from_skid_rdy | __axi_reader__axi_st_s_data_has_been_sent_reg) & (~p1_and_1929 | axi_reader__resp_s_data_from_skid_rdy | __axi_reader__resp_s_data_has_been_sent_reg);
  assign and_2094 = ((and_2070 | 16'h0200) & {16{p0_____state_4__1 < 4'ha}} | 16'h0400) & {16{p0_____state_4__1 < 4'hb}};
  assign p2_stage_done = p1_valid & or_2416 & p2_all_active_outputs_ready;
  assign p2_not_valid = ~p1_valid;
  assign is_last_group = ____state_3 == 8'h00;
  assign not_1927 = ~____state_0;
  assign p1_enable = p2_stage_done | p2_not_valid;
  assign and_1929 = ____state_0 & is_last_group;
  assign nor_1930 = ~(not_1927 | is_last_group);
  assign sel_1900 = ____state_5 > 4'h2 ? 3'h7 : {1'h0, |____state_5[3:1] ? 2'h3 : {1'h0, ____state_5 != 4'h0}};
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign concat_2156 = {1'h0, p1_ugt_2110 ? 13'h1fff : {1'h0, p1_ugt_2102 ? 12'hfff : {1'h0, p1_sel_2098}}};
  assign ____state_2__next_value_predicates = {not_1927, and_1929};
  assign ____state_3__next_value_predicates = {not_1927, nor_1930, and_1929};
  assign ____state_4__next_value_predicates = {not_1927, ____state_0};
  assign concat_2068 = {1'h0, p0_____state_5__1[3] ? 8'hff : {1'h0, p0_ugt_1918 ? 7'h7f : {1'h0, p0_sel_1917}}};
  assign MAX_LANE__2 = 4'hf;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_stage_done = ____state_0 | __axi_reader__conf_r_data_valid_reg | __axi_reader__conf_r_data_valid_skid_reg;
  assign one_hot_1937 = {____state_2__next_value_predicates[1:0] == 2'h0, ____state_2__next_value_predicates[1] && !____state_2__next_value_predicates[0], ____state_2__next_value_predicates[0]};
  assign one_hot_1938 = {____state_3__next_value_predicates[2:0] == 3'h0, ____state_3__next_value_predicates[2] && ____state_3__next_value_predicates[1:0] == 2'h0, ____state_3__next_value_predicates[1] && !____state_3__next_value_predicates[0], ____state_3__next_value_predicates[0]};
  assign one_hot_1939 = {____state_4__next_value_predicates[1:0] == 2'h0, ____state_4__next_value_predicates[1] && !____state_4__next_value_predicates[0], ____state_4__next_value_predicates[0]};
  assign and_2111 = ((and_2094 | 16'h0800) & {16{p0_____state_4__1 < 4'hc}} | 16'h1000) & {16{p0_____state_4__1 < 4'hd}};
  assign p0_data_enable = p0_enable & p0_stage_done;
  assign __axi_reader__axi_st_s_vld_buf = or_2416 & p1_valid & nor_2181;
  assign __axi_reader__axi_st_s_data_not_has_been_sent = ~__axi_reader__axi_st_s_data_has_been_sent_reg;
  assign __axi_reader__resp_s_vld_buf = or_2416 & p1_valid & p1_and_1929;
  assign __axi_reader__resp_s_data_not_has_been_sent = ~__axi_reader__resp_s_data_has_been_sent_reg;
  assign axi_reader__conf_r_data_select = __axi_reader__conf_r_data_valid_skid_reg ? __axi_reader__conf_r_data_skid_reg : __axi_reader__conf_r_data_reg;
  assign axi_reader__conf_r_data_from_skid_rdy = ~__axi_reader__conf_r_data_valid_skid_reg;
  assign and_2270 = not_1927 & p0_data_enable;
  assign axi_reader__axi_r_r_data_from_skid_rdy = ~__axi_reader__axi_r_r_data_valid_skid_reg;
  assign and_2271 = p1_____state_0__1 & p2_stage_done;
  assign high_mask_squeezed = p1_eq_1928 ? 15'h7fff : {1'h0, p1_ugt_2118 ? 14'h3fff : concat_2156};
  assign high_mask_squeezed_const_lsb_bits = 1'h1;
  assign __axi_reader__axi_st_s_data_valid_and_not_has_been_sent = __axi_reader__axi_st_s_vld_buf & __axi_reader__axi_st_s_data_not_has_been_sent;
  assign __axi_reader__resp_s_data_valid_and_not_has_been_sent = __axi_reader__resp_s_vld_buf & __axi_reader__resp_s_data_not_has_been_sent;
  assign MAX_LANE = 4'hf;
  assign and_2242 = and_1929 & p0_data_enable;
  assign axi_reader__conf_r_select = not_1927 ? axi_reader__conf_r_data_select : literal_1942;
  assign and_2249 = nor_1930 & p0_data_enable;
  assign and_2256 = ____state_0 & p0_data_enable;
  assign axi_reader__conf_r_data_data_valid_load_en = axi_reader__conf_r_vld & axi_reader__conf_r_data_from_skid_rdy;
  assign axi_reader__conf_r_data_to_is_not_rdy = ~and_2270;
  assign axi_reader__axi_r_r_data_data_valid_load_en = axi_reader__axi_r_r_vld & axi_reader__axi_r_r_data_from_skid_rdy;
  assign axi_reader__axi_r_r_data_to_is_not_rdy = ~and_2271;
  assign low_mask = p1_and_2124 | 16'h8000;
  assign high_mask = {high_mask_squeezed, high_mask_squeezed_const_lsb_bits};
  assign axi_reader__axi_st_s_data_data_valid_load_en = __axi_reader__axi_st_s_data_valid_and_not_has_been_sent & axi_reader__axi_st_s_data_from_skid_rdy;
  assign axi_reader__axi_st_s_data_to_is_not_rdy = ~axi_reader__axi_st_s_rdy;
  assign axi_reader__resp_s_data_data_valid_load_en = __axi_reader__resp_s_data_valid_and_not_has_been_sent & axi_reader__resp_s_data_from_skid_rdy;
  assign axi_reader__resp_s_data_to_is_not_rdy = ~axi_reader__resp_s_rdy;
  assign ____state_2__at_most_one_next_value = not_1927 == one_hot_1937[1] & and_1929 == one_hot_1937[0];
  assign ____state_3__at_most_one_next_value = not_1927 == one_hot_1938[2] & nor_1930 == one_hot_1938[1] & and_1929 == one_hot_1938[0];
  assign ____state_4__at_most_one_next_value = not_1927 == one_hot_1939[1] & ____state_0 == one_hot_1939[0];
  assign concat_2092 = {1'h0, p0_____state_5__1 > 4'h9 ? 10'h3ff : {1'h0, p0_____state_5__1 > 4'h8 ? 9'h1ff : concat_2068}};
  assign concat_1914 = {1'h0, ____state_5 > 4'h4 ? 5'h1f : {1'h0, |____state_5[3:2] ? MAX_LANE__2 : {1'h0, sel_1900}}};
  assign high_lane = is_last_group ? ____state_5 : MAX_LANE;
  assign MAX_LANE__1 = 4'hf;
  assign is_last_tran = ____state_2 == 16'h0000;
  assign concat_2244 = {and_2270, and_2242};
  assign concat_2251 = {and_2270, and_2249, and_2242};
  assign add_1968 = ____state_3 + 8'hff;
  assign concat_2257 = {and_2270, and_2256};
  assign __axi_reader__axi_st_s_data_valid_and_all_active_outputs_ready = __axi_reader__axi_st_s_vld_buf & p2_all_active_outputs_ready;
  assign __axi_reader__resp_s_data_valid_and_all_active_outputs_ready = __axi_reader__resp_s_vld_buf & p2_all_active_outputs_ready;
  assign axi_reader__conf_r_data_data_is_sent_to = __axi_reader__conf_r_data_valid_reg & and_2270 & axi_reader__conf_r_data_from_skid_rdy;
  assign axi_reader__conf_r_data_skid_data_load_en = __axi_reader__conf_r_data_valid_reg & axi_reader__conf_r_data_data_valid_load_en & axi_reader__conf_r_data_to_is_not_rdy;
  assign axi_reader__conf_r_data_skid_valid_set_zero = __axi_reader__conf_r_data_valid_skid_reg & and_2270;
  assign axi_reader__axi_r_r_data_data_is_sent_to = __axi_reader__axi_r_r_data_valid_reg & and_2271 & axi_reader__axi_r_r_data_from_skid_rdy;
  assign axi_reader__axi_r_r_data_skid_data_load_en = __axi_reader__axi_r_r_data_valid_reg & axi_reader__axi_r_r_data_data_valid_load_en & axi_reader__axi_r_r_data_to_is_not_rdy;
  assign axi_reader__axi_r_r_data_skid_valid_set_zero = __axi_reader__axi_r_r_data_valid_skid_reg & and_2271;
  assign axi_r_data = axi_reader__axi_r_r_select[131:4];
  assign mask = low_mask & high_mask;
  assign axi_reader__axi_st_s_data_data_is_sent_to = __axi_reader__axi_st_s_data_valid_reg & axi_reader__axi_st_s_rdy & axi_reader__axi_st_s_data_from_skid_rdy;
  assign axi_reader__axi_st_s_data_skid_data_load_en = __axi_reader__axi_st_s_data_valid_reg & axi_reader__axi_st_s_data_data_valid_load_en & axi_reader__axi_st_s_data_to_is_not_rdy;
  assign axi_reader__axi_st_s_data_skid_valid_set_zero = __axi_reader__axi_st_s_data_valid_skid_reg & axi_reader__axi_st_s_rdy;
  assign axi_reader__resp_s_data_data_is_sent_to = __axi_reader__resp_s_data_valid_reg & axi_reader__resp_s_rdy & axi_reader__resp_s_data_from_skid_rdy;
  assign axi_reader__resp_s_data_skid_data_load_en = __axi_reader__resp_s_data_valid_reg & axi_reader__resp_s_data_data_valid_load_en & axi_reader__resp_s_data_to_is_not_rdy;
  assign axi_reader__resp_s_data_skid_valid_set_zero = __axi_reader__resp_s_data_valid_skid_reg & axi_reader__resp_s_rdy;
  assign axi_reader__axi_st_s_data_select = __axi_reader__axi_st_s_data_valid_skid_reg ? __axi_reader__axi_st_s_data_skid_reg : __axi_reader__axi_st_s_data_reg;
  assign axi_reader__axi_st_s_data_valid_or = __axi_reader__axi_st_s_data_valid_reg | __axi_reader__axi_st_s_data_valid_skid_reg;
  assign axi_reader__resp_s_data_select = __axi_reader__resp_s_data_valid_skid_reg ? __axi_reader__resp_s_data_skid_reg : __axi_reader__resp_s_data_reg;
  assign axi_reader__resp_s_data_valid_or = __axi_reader__resp_s_data_valid_reg | __axi_reader__resp_s_data_valid_skid_reg;
  assign or_2408 = ~p0_stage_done | ____state_2__at_most_one_next_value | rst;
  assign sel_2098 = p0_____state_5__1 > 4'ha ? 11'h7ff : concat_2092;
  assign ugt_2102 = p0_____state_5__1 > 4'hb;
  assign ugt_2110 = p0_____state_5__1 > 4'hc;
  assign ugt_2118 = p0_____state_5__1 > 4'hd;
  assign and_2124 = ((and_2111 | 16'h2000) & {16{p0_____state_4__1 < 4'he}} | 16'h4000) & {16{~(&p0_____state_4__1)}};
  assign eq_1885 = ____state_4[3:1] == 3'h0;
  assign sel_1917 = ____state_5 > 4'h5 ? 6'h3f : concat_1914;
  assign ugt_1918 = ____state_5 > 4'h6;
  assign eq_1928 = high_lane == MAX_LANE__1;
  assign and_1940 = is_last_group & is_last_tran;
  assign nand_1961 = ~(____state_0 & is_last_group);
  assign one_hot_sel_2245 = 16'h0000 & {16{concat_2244[0]}} | axi_reader__conf_r_select[31:16] & {16{concat_2244[1]}};
  assign or_2246 = and_2270 | and_2242;
  assign one_hot_sel_2252 = 8'h00 & {8{concat_2251[0]}} | add_1968 & {8{concat_2251[1]}} | axi_reader__conf_r_select[15:8] & {8{concat_2251[2]}};
  assign or_2253 = and_2270 | and_2249 | and_2242;
  assign one_hot_sel_2258 = 4'h0 & {4{concat_2257[0]}} | axi_reader__conf_r_select[7:4] & {4{concat_2257[1]}};
  assign or_2259 = and_2270 | and_2256;
  assign one_hot_sel_2265 = 4'h0 & {4{concat_2244[0]}} | axi_reader__conf_r_select[3:0] & {4{concat_2244[1]}};
  assign __axi_reader__axi_st_s_data_not_stage_load = ~__axi_reader__axi_st_s_data_valid_and_all_active_outputs_ready;
  assign __axi_reader__axi_st_s_data_has_been_sent_reg_load_en = axi_reader__axi_st_s_data_data_valid_load_en | __axi_reader__axi_st_s_data_valid_and_all_active_outputs_ready;
  assign __axi_reader__resp_s_data_not_stage_load = ~__axi_reader__resp_s_data_valid_and_all_active_outputs_ready;
  assign __axi_reader__resp_s_data_has_been_sent_reg_load_en = axi_reader__resp_s_data_data_valid_load_en | __axi_reader__resp_s_data_valid_and_all_active_outputs_ready;
  assign axi_reader__conf_r_data_data_valid_load_en__1 = axi_reader__conf_r_data_data_is_sent_to | axi_reader__conf_r_data_data_valid_load_en;
  assign axi_reader__conf_r_data_skid_valid_load_en = axi_reader__conf_r_data_skid_data_load_en | axi_reader__conf_r_data_skid_valid_set_zero;
  assign axi_reader__axi_r_r_data_data_valid_load_en__1 = axi_reader__axi_r_r_data_data_is_sent_to | axi_reader__axi_r_r_data_data_valid_load_en;
  assign axi_reader__axi_r_r_data_skid_valid_load_en = axi_reader__axi_r_r_data_skid_data_load_en | axi_reader__axi_r_r_data_skid_valid_set_zero;
  assign __axi_reader__axi_st_s_data_buf = {axi_r_data, mask, mask, 8'h00, 8'h00, p1_and_1940};
  assign axi_reader__axi_st_s_data_data_valid_load_en__1 = axi_reader__axi_st_s_data_data_is_sent_to | axi_reader__axi_st_s_data_data_valid_load_en;
  assign axi_reader__axi_st_s_data_skid_valid_load_en = axi_reader__axi_st_s_data_skid_data_load_en | axi_reader__axi_st_s_data_skid_valid_set_zero;
  assign axi_reader__resp_s_data_data_valid_load_en__1 = axi_reader__resp_s_data_data_is_sent_to | axi_reader__resp_s_data_data_valid_load_en;
  assign axi_reader__resp_s_data_skid_valid_load_en = axi_reader__resp_s_data_skid_data_load_en | axi_reader__resp_s_data_skid_valid_set_zero;
  always @ (posedge clk) begin
    if (rst) begin
      ____state_4 <= 4'h0;
      ____state_5 <= 4'h0;
      ____state_3 <= 8'h00;
      ____state_0 <= 1'h0;
      ____state_2 <= 16'h0000;
      p0_____state_0__1 <= 1'h0;
      p0_____state_4__1 <= 4'h0;
      p0_____state_5__1 <= 4'h0;
      p0_eq_1885 <= 1'h0;
      p0_sel_1917 <= 6'h00;
      p0_ugt_1918 <= 1'h0;
      p0_eq_1928 <= 1'h0;
      p0_not_1927 <= 1'h0;
      p0_and_1940 <= 1'h0;
      p0_and_1929 <= 1'h0;
      p1_____state_0__1 <= 1'h0;
      p1_sel_2098 <= 11'h000;
      p1_ugt_2102 <= 1'h0;
      p1_ugt_2110 <= 1'h0;
      p1_ugt_2118 <= 1'h0;
      p1_eq_1928 <= 1'h0;
      p1_and_2124 <= 16'h0000;
      p1_not_1927 <= 1'h0;
      p1_and_1940 <= 1'h0;
      p1_and_1929 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      __axi_reader__axi_st_s_data_has_been_sent_reg <= 1'h0;
      __axi_reader__resp_s_data_has_been_sent_reg <= 1'h0;
      __axi_reader__conf_r_data_reg <= __axi_reader__conf_r_data_reg_init;
      __axi_reader__conf_r_data_skid_reg <= __axi_reader__conf_r_data_skid_reg_init;
      __axi_reader__conf_r_data_valid_reg <= 1'h0;
      __axi_reader__conf_r_data_valid_skid_reg <= 1'h0;
      __axi_reader__axi_r_r_data_reg <= __axi_reader__axi_r_r_data_reg_init;
      __axi_reader__axi_r_r_data_skid_reg <= __axi_reader__axi_r_r_data_skid_reg_init;
      __axi_reader__axi_r_r_data_valid_reg <= 1'h0;
      __axi_reader__axi_r_r_data_valid_skid_reg <= 1'h0;
      __axi_reader__axi_st_s_data_reg <= __axi_reader__axi_st_s_data_reg_init;
      __axi_reader__axi_st_s_data_skid_reg <= __axi_reader__axi_st_s_data_skid_reg_init;
      __axi_reader__axi_st_s_data_valid_reg <= 1'h0;
      __axi_reader__axi_st_s_data_valid_skid_reg <= 1'h0;
      __axi_reader__resp_s_data_reg <= 1'h0;
      __axi_reader__resp_s_data_skid_reg <= 1'h0;
      __axi_reader__resp_s_data_valid_reg <= 1'h0;
      __axi_reader__resp_s_data_valid_skid_reg <= 1'h0;
    end else begin
      ____state_4 <= or_2259 ? one_hot_sel_2258 : ____state_4;
      ____state_5 <= or_2246 ? one_hot_sel_2265 : ____state_5;
      ____state_3 <= or_2253 ? one_hot_sel_2252 : ____state_3;
      ____state_0 <= p0_data_enable ? nand_1961 : ____state_0;
      ____state_2 <= or_2246 ? one_hot_sel_2245 : ____state_2;
      p0_____state_0__1 <= p0_data_enable ? ____state_0 : p0_____state_0__1;
      p0_____state_4__1 <= p0_data_enable ? ____state_4 : p0_____state_4__1;
      p0_____state_5__1 <= p0_data_enable ? ____state_5 : p0_____state_5__1;
      p0_eq_1885 <= p0_data_enable ? eq_1885 : p0_eq_1885;
      p0_sel_1917 <= p0_data_enable ? sel_1917 : p0_sel_1917;
      p0_ugt_1918 <= p0_data_enable ? ugt_1918 : p0_ugt_1918;
      p0_eq_1928 <= p0_data_enable ? eq_1928 : p0_eq_1928;
      p0_not_1927 <= p0_data_enable ? not_1927 : p0_not_1927;
      p0_and_1940 <= p0_data_enable ? and_1940 : p0_and_1940;
      p0_and_1929 <= p0_data_enable ? and_1929 : p0_and_1929;
      p1_____state_0__1 <= p1_data_enable ? p0_____state_0__1 : p1_____state_0__1;
      p1_sel_2098 <= p1_data_enable ? sel_2098 : p1_sel_2098;
      p1_ugt_2102 <= p1_data_enable ? ugt_2102 : p1_ugt_2102;
      p1_ugt_2110 <= p1_data_enable ? ugt_2110 : p1_ugt_2110;
      p1_ugt_2118 <= p1_data_enable ? ugt_2118 : p1_ugt_2118;
      p1_eq_1928 <= p1_data_enable ? p0_eq_1928 : p1_eq_1928;
      p1_and_2124 <= p1_data_enable ? and_2124 : p1_and_2124;
      p1_not_1927 <= p1_data_enable ? p0_not_1927 : p1_not_1927;
      p1_and_1940 <= p1_data_enable ? p0_and_1940 : p1_and_1940;
      p1_and_1929 <= p1_data_enable ? p0_and_1929 : p1_and_1929;
      p0_valid <= p0_enable ? p0_stage_done : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      __axi_reader__axi_st_s_data_has_been_sent_reg <= __axi_reader__axi_st_s_data_has_been_sent_reg_load_en ? __axi_reader__axi_st_s_data_not_stage_load : __axi_reader__axi_st_s_data_has_been_sent_reg;
      __axi_reader__resp_s_data_has_been_sent_reg <= __axi_reader__resp_s_data_has_been_sent_reg_load_en ? __axi_reader__resp_s_data_not_stage_load : __axi_reader__resp_s_data_has_been_sent_reg;
      __axi_reader__conf_r_data_reg <= axi_reader__conf_r_data_data_valid_load_en ? axi_reader__conf_r_data : __axi_reader__conf_r_data_reg;
      __axi_reader__conf_r_data_skid_reg <= axi_reader__conf_r_data_skid_data_load_en ? __axi_reader__conf_r_data_reg : __axi_reader__conf_r_data_skid_reg;
      __axi_reader__conf_r_data_valid_reg <= axi_reader__conf_r_data_data_valid_load_en__1 ? axi_reader__conf_r_vld : __axi_reader__conf_r_data_valid_reg;
      __axi_reader__conf_r_data_valid_skid_reg <= axi_reader__conf_r_data_skid_valid_load_en ? axi_reader__conf_r_data_from_skid_rdy : __axi_reader__conf_r_data_valid_skid_reg;
      __axi_reader__axi_r_r_data_reg <= axi_reader__axi_r_r_data_data_valid_load_en ? axi_reader__axi_r_r_data : __axi_reader__axi_r_r_data_reg;
      __axi_reader__axi_r_r_data_skid_reg <= axi_reader__axi_r_r_data_skid_data_load_en ? __axi_reader__axi_r_r_data_reg : __axi_reader__axi_r_r_data_skid_reg;
      __axi_reader__axi_r_r_data_valid_reg <= axi_reader__axi_r_r_data_data_valid_load_en__1 ? axi_reader__axi_r_r_vld : __axi_reader__axi_r_r_data_valid_reg;
      __axi_reader__axi_r_r_data_valid_skid_reg <= axi_reader__axi_r_r_data_skid_valid_load_en ? axi_reader__axi_r_r_data_from_skid_rdy : __axi_reader__axi_r_r_data_valid_skid_reg;
      __axi_reader__axi_st_s_data_reg <= axi_reader__axi_st_s_data_data_valid_load_en ? __axi_reader__axi_st_s_data_buf : __axi_reader__axi_st_s_data_reg;
      __axi_reader__axi_st_s_data_skid_reg <= axi_reader__axi_st_s_data_skid_data_load_en ? __axi_reader__axi_st_s_data_reg : __axi_reader__axi_st_s_data_skid_reg;
      __axi_reader__axi_st_s_data_valid_reg <= axi_reader__axi_st_s_data_data_valid_load_en__1 ? __axi_reader__axi_st_s_data_valid_and_not_has_been_sent : __axi_reader__axi_st_s_data_valid_reg;
      __axi_reader__axi_st_s_data_valid_skid_reg <= axi_reader__axi_st_s_data_skid_valid_load_en ? axi_reader__axi_st_s_data_from_skid_rdy : __axi_reader__axi_st_s_data_valid_skid_reg;
      __axi_reader__resp_s_data_reg <= axi_reader__resp_s_data_data_valid_load_en ? is_err : __axi_reader__resp_s_data_reg;
      __axi_reader__resp_s_data_skid_reg <= axi_reader__resp_s_data_skid_data_load_en ? __axi_reader__resp_s_data_reg : __axi_reader__resp_s_data_skid_reg;
      __axi_reader__resp_s_data_valid_reg <= axi_reader__resp_s_data_data_valid_load_en__1 ? __axi_reader__resp_s_data_valid_and_not_has_been_sent : __axi_reader__resp_s_data_valid_reg;
      __axi_reader__resp_s_data_valid_skid_reg <= axi_reader__resp_s_data_skid_valid_load_en ? axi_reader__resp_s_data_from_skid_rdy : __axi_reader__resp_s_data_valid_skid_reg;
    end
  end
  assign axi_reader__axi_r_r_rdy = axi_reader__axi_r_r_data_from_skid_rdy;
  assign axi_reader__axi_st_s_data = axi_reader__axi_st_s_data_select;
  assign axi_reader__axi_st_s_vld = axi_reader__axi_st_s_data_valid_or;
  assign axi_reader__conf_r_rdy = axi_reader__conf_r_data_from_skid_rdy;
  assign axi_reader__resp_s_data = axi_reader__resp_s_data_select;
  assign axi_reader__resp_s_vld = axi_reader__resp_s_data_valid_or;
endmodule


module __xls_modules_zstd_memory_axi_reader__MemReaderAdvNoFsmInst__MemReaderAdvNoFsm_0__AxiReaderNoFsm_0__AxiReaderInternalR_0__16_128_16_8_8_5_4_12_next(
  input wire clk,
  input wire rst,
  input wire [139:0] mem_reader__axi_r_r_data,
  input wire mem_reader__axi_r_r_vld,
  input wire mem_reader__axi_st_in_rdy,
  input wire [47:0] mem_reader__rconf_data,
  input wire mem_reader__rconf_vld,
  input wire mem_reader__rresp_rdy,
  output wire mem_reader__axi_r_r_rdy,
  output wire [176:0] mem_reader__axi_st_in_data,
  output wire mem_reader__axi_st_in_vld,
  output wire mem_reader__rconf_rdy,
  output wire mem_reader__rresp_data,
  output wire mem_reader__rresp_vld
);
  // ===== Instantiations
  __axi_reader__AxiReaderInternalRInst__AxiReaderInternalR_0__16_128_16_8_8_5_4_12_next __axi_reader__AxiReaderInternalRInst__AxiReaderInternalR_0__16_128_16_8_8_5_4_12_next_inst0 (
    .rst(rst),
    .axi_reader__axi_r_r_data(mem_reader__axi_r_r_data),
    .axi_reader__axi_r_r_vld(mem_reader__axi_r_r_vld),
    .axi_reader__axi_st_s_rdy(mem_reader__axi_st_in_rdy),
    .axi_reader__conf_r_data(mem_reader__rconf_data),
    .axi_reader__conf_r_vld(mem_reader__rconf_vld),
    .axi_reader__resp_s_rdy(mem_reader__rresp_rdy),
    .axi_reader__axi_r_r_rdy(mem_reader__axi_r_r_rdy),
    .axi_reader__axi_st_s_data(mem_reader__axi_st_in_data),
    .axi_reader__axi_st_s_vld(mem_reader__axi_st_in_vld),
    .axi_reader__conf_r_rdy(mem_reader__rconf_rdy),
    .axi_reader__resp_s_data(mem_reader__rresp_data),
    .axi_reader__resp_s_vld(mem_reader__rresp_vld),
    .clk(clk)
  );

endmodule
